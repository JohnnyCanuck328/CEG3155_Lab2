library verilog;
use verilog.vl_types.all;
entity eightBitAddSub_vlg_vec_tst is
end eightBitAddSub_vlg_vec_tst;
