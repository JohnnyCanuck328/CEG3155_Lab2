library verilog;
use verilog.vl_types.all;
entity twoComp_vlg_vec_tst is
end twoComp_vlg_vec_tst;
