library verilog;
use verilog.vl_types.all;
entity divider4bit_vlg_vec_tst is
end divider4bit_vlg_vec_tst;
