library verilog;
use verilog.vl_types.all;
entity twoComp_vlg_sample_tst is
    port(
        A               : in     vl_logic_vector(3 downto 0);
        enable          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end twoComp_vlg_sample_tst;
