library verilog;
use verilog.vl_types.all;
entity fullSubtractor_vlg_check_tst is
    port(
        Bout            : in     vl_logic;
        D               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end fullSubtractor_vlg_check_tst;
