library verilog;
use verilog.vl_types.all;
entity multiplier4bit_vlg_vec_tst is
end multiplier4bit_vlg_vec_tst;
