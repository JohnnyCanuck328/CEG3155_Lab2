library verilog;
use verilog.vl_types.all;
entity fourBitMulti_vlg_vec_tst is
end fourBitMulti_vlg_vec_tst;
