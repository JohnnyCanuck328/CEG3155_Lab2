library verilog;
use verilog.vl_types.all;
entity fourBitMulti_vlg_check_tst is
    port(
        product         : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end fourBitMulti_vlg_check_tst;
