library verilog;
use verilog.vl_types.all;
entity eightbitaddsub_vlg_vec_tst is
end eightbitaddsub_vlg_vec_tst;
