library verilog;
use verilog.vl_types.all;
entity divider4bit_vlg_check_tst is
    port(
        quotient        : in     vl_logic_vector(3 downto 0);
        remainder       : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end divider4bit_vlg_check_tst;
