library verilog;
use verilog.vl_types.all;
entity fullSubtractor_vlg_vec_tst is
end fullSubtractor_vlg_vec_tst;
