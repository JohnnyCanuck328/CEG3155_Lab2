library verilog;
use verilog.vl_types.all;
entity fourbitaddsub_vlg_vec_tst is
end fourbitaddsub_vlg_vec_tst;
