library verilog;
use verilog.vl_types.all;
entity twoAnd_vlg_vec_tst is
end twoAnd_vlg_vec_tst;
