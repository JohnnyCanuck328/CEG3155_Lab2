library verilog;
use verilog.vl_types.all;
entity multiplier4bit_vlg_check_tst is
    port(
        P               : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end multiplier4bit_vlg_check_tst;
