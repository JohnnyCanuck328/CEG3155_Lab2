library verilog;
use verilog.vl_types.all;
entity twoComp8bit_vlg_vec_tst is
end twoComp8bit_vlg_vec_tst;
